LIBRARY ieee;
USE ieee.std_logic_1164.all;
-- Simple module that connects the SW switches to the LEDR lights

ENTITY PLab1_Parte1 IS

PORT ( SW : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
LEDR : OUT STD_LOGIC_VECTOR(17 DOWNTO 0)); -- red LEDs
END ;
ARCHITECTURE Behavior OF PLab1_Parte1 IS
BEGIN
LEDR <= SW;
END Behavior;